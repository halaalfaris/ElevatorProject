//4-1 Mux

module mux1 (i0,i1,i2,i3,s0,s1,out);
input i0,i1,i2,i3,s0,s1;
output out;
 assign out = i0&~s0&~s1 |i1&s0&~s1 |i2&~s0&s1 |i3&s0&s1;

endmodule